class sr_monitor extends uvm_monitor; 

  //---------------------------------------------------------------------------- 

  `uvm_component_utils(sr_monitor) 

  //---------------------------------------------------------------------------- 

 

  //------------------- constructor -------------------------------------------- 

  function new(string name="sr_monitor",uvm_component parent); 

    super.new(name,parent); 

  endfunction 

  //---------------------------------------------------------------------------- 

   

  //---------------- sequence_item class --------------------------------------- 

  sr_sequence_item  txn; 

  //---------------------------------------------------------------------------- 

   

  //------------------------ virtual interface handle---------------------------   

  virtual interface intf vif; 

  //---------------------------------------------------------------------------- 

 

  //------------------------ analysis port ------------------------------------- 

  uvm_analysis_port#(sr_sequence_item) ap_mon; 

  //---------------------------------------------------------------------------- 

   

  //------------------- build phase -------------------------------------------- 

  function void build_phase(uvm_phase phase); 

    super.build_phase(phase); 

    if(!(uvm_config_db#(virtual intf)::get(this,"","vif",vif))) 

    begin 

      `uvm_fatal("monitor","unable to get interface") 

    end 

     

    ap_mon=new("ap_mon",this); 

  endfunction 

  //---------------------------------------------------------------------------- 

 

  //-------------------- run phase --------------------------------------------- 

  task run_phase(uvm_phase phase); 

    sr_sequence_item txn=sr_sequence_item::type_id::create("txn"); 

    forever 

    begin 

      sample_dut(txn); 

      ap_mon.write(txn); 

    end 

  endtask 

  //---------------------------------------------------------------------------- 

 

  task sample_dut(output sr_sequence_item txn); 

    sr_sequence_item t = sr_sequence_item::type_id::create("t"); 

    #5.1; 

    t.s    = vif.s; 

    t.r    = vif.r; 

    t.q    = vif.q; 

    t.qbar = vif.qbar; 

    txn    = t; 

  endtask : sample_dut 

 

endclass:sr_monitor 
